//29-6

`include "interface.sv"
`include "random_test.sv"

module tb_top;
  
  bit rdclk;
  bit wrclk;
  bit wrst_n, rrst_n;
//   bit wr_en, rd_en;

  //Clock signals
  
  
  
  //Reset Signals
  initial begin
    rdclk=1'b0;
    wrclk=1'b0;
    wrst_n=1'b0;
    rrst_n=1'b0;
    #30 wrst_n=1'b1;
    rrst_n=1'b1;
//     #40 wrst_n=1'b0; 
//     #5 rrst_n=1'b0;
//      #10 wrst_n=1'b1;
//     #5 rrst_n=1'b1;
  end
  
  always begin  #25 rdclk= ~rdclk; end     
  always begin  #10 wrclk= ~wrclk; end

  //Enable Signals
  //initial begin
//     #35 rd_en=1'b1; wr_en=1'b0;
//     #35 rd_en=1'b0; wr_en=1'b1;
//     #35 rd_en=1'b1; wr_en=1'b0;
//     #35 rd_en=1'b0; wr_en=1'b1;
//     #35 rd_en=1'b1; wr_en=1'b0;
//     #35 rd_en=1'b0; wr_en=1'b1;
//     #35 rd_en=1'b1; wr_en=1'b0;
//     #35 rd_en=1'b0; wr_en=1'b1;
//     #35 rd_en=1'b1; wr_en=1'b0;
    
//      #40 wr_en=1'b1;
//     #60 rd_en = 1'b1; 
    
  //end

  
  fifo_intf vif(wrclk,rdclk,wrst_n,rrst_n);
  test t1(vif);
  
  asynchronous_fifo fifo_instance  (
    .wrclk(vif.wrclk),
    .rdclk(vif.rdclk),
    .wrst_n(vif.wrst_n),
    .rrst_n(vif.rrst_n),
    .wr_en(vif.wr_en),
    .rd_en(vif.rd_en),
    .data_in(vif.data_in),
    .data_out(vif.data_out),
    .fifo_full(vif.fifo_full),
    .fifo_empty(vif.fifo_empty)
  );
  
  
  initial begin 
    $dumpfile("dump.vcd");
    $dumpvars;
  end
 
endmodule